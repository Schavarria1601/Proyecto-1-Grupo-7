`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/02/2017 04:20:05 PM
// Design Name: 
// Module Name: Font_Rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module font_rom(
    clk,
    addr,
    rom_data
    );
    
    //  Parametrizacion del bus de datos.
    parameter bus_addr = 7;     //  OJO, aqui puede que exista un problema.
    parameter bus_data = 32;
    //  Declaracion de entradas y salidas.
    input wire clk;
    input wire [bus_addr-1:0] addr;
    output reg [bus_data-1:0] rom_data;
    
    //Número de fila seleccionado por rom_addr
    reg [bus_addr-1:0] addr_reg;
    
    always @(posedge clk)
        addr_reg <= addr;
        
    always @*
            case(addr_reg)
                7'h00: rom_data = 32'b01111111111111111111111111000000;
                7'h01: rom_data = 32'b01111111111111111111111111000000;
                7'h02: rom_data = 32'b01111111111111111111111111000000;
                7'h03: rom_data = 32'b01111111111111111111111111000000;
                7'h04: rom_data = 32'b01111100000000000111111111111000;
                7'h05: rom_data = 32'b01111100000000000111111111111000;
                7'h06: rom_data = 32'b01111100000000000111111111111000;
                7'h07: rom_data = 32'b01111100000000000111111111111000;
                7'h08: rom_data = 32'b01111100000000000111111111111000;
                7'h09: rom_data = 32'b01111100000000000111111111111000; 
                7'h0A: rom_data = 32'b01111100000000000111111111111000;
                7'h0B: rom_data = 32'b01111100000000000111111111111000;
                7'h0C: rom_data = 32'b01111100000000000111111111111000;
                7'h0D: rom_data = 32'b01111100000000000111111111111000;
                7'h0E: rom_data = 32'b01111100000000000111111111111000;
                7'h0F: rom_data = 32'b01111100000000000111111111111000;
                7'h10: rom_data = 32'b01111100000000000111111111111000;
                7'h11: rom_data = 32'b01111100000000000111111111111000;
                7'h12: rom_data = 32'b01111100000000000111111111111000;
                7'h13: rom_data = 32'b01111100000000000111111111111000;
                7'h14: rom_data = 32'b01111100000000000111111111111000;
                7'h15: rom_data = 32'b01111100000000000111111111111000;
                7'h16: rom_data = 32'b01111100000000000111111111111000;
                7'h17: rom_data = 32'b01111100000000000111111111111000;
                7'h18: rom_data = 32'b01111100000000000111111111111000;
                7'h19: rom_data = 32'b01111100000000000111111111111000;
                7'h1a: rom_data = 32'b01111100000000000111111111111000;
                7'h1b: rom_data = 32'b01111100000000000111111111111000;
                7'h1c: rom_data = 32'b01111111111111111111111111000000;
                7'h1d: rom_data = 32'b01111111111111111111111111000000;
                7'h1e: rom_data = 32'b01111111111111111111111111000000;
                7'h1f: rom_data = 32'b00000000000000000000000000000000;
            
            
                7'h20: rom_data = 32'b00011111111111111111111111110000;
                7'h21: rom_data = 32'b00011111111111111111111111110000;
                7'h22: rom_data = 32'b00011111111111111111111111110000;
                7'h23: rom_data = 32'b01111111111111111111111111110000;
                7'h24: rom_data = 32'b01111100000000000000000000000000;
                7'h25: rom_data = 32'b01111100000000000000000000000000;
                7'h26: rom_data = 32'b01111100000000000000000000000000;
                7'h27: rom_data = 32'b01111100000000000000000000000000;
                7'h28: rom_data = 32'b01111100000000000000000000000000;
                7'h29: rom_data = 32'b01111100000000000000000000000000; 
                7'h2a: rom_data = 32'b01111100000000000000000000000000;
                7'h2b: rom_data = 32'b01111100011111111111111111111000;
                7'h2c: rom_data = 32'b01111100011111111111111111111000;
                7'h2d: rom_data = 32'b01111100011111111111111111111000;
                7'h2e: rom_data = 32'b01111100011111111111111111111000;
                7'h2f: rom_data = 32'b01111100011111111111111111111000;
                7'h30: rom_data = 32'b01111100000000000111111111111000;
                7'h31: rom_data = 32'b01111100000000000111111111111000;
                7'h32: rom_data = 32'b01111100000000000111111111111000;
                7'h33: rom_data = 32'b01111100000000000111111111111000;
                7'h34: rom_data = 32'b01111100000000000111111111111000;
                7'h35: rom_data = 32'b01111100000000000111111111111000;
                7'h36: rom_data = 32'b01111100000000000111111111111000;
                7'h37: rom_data = 32'b01111100000000000111111111111000;
                7'h38: rom_data = 32'b01111100000000000111111111111000;
                7'h39: rom_data = 32'b01111100000000000111111111111000;
                7'h3a: rom_data = 32'b01111100000000000111111111111000;
                7'h3b: rom_data = 32'b01111111111111111111111111111000;
                7'h3c: rom_data = 32'b01111111111111111111111111111000;
                7'h3d: rom_data = 32'b00011111111111111111111111111000;
                7'h3e: rom_data = 32'b00011111111111111111111111111000;
                7'h3f: rom_data = 32'b00000000000000000000000000000000;
                
              
                7'h40: rom_data = 32'b00001111111111111111111111111111;
                7'h41: rom_data = 32'b00001111111111111111111111111111;
                7'h42: rom_data = 32'b01111111111111111111111111111111;
                7'h43: rom_data = 32'b01111111111111111111111111111111;
                7'h44: rom_data = 32'b01111111111111111111111111111111;
                7'h45: rom_data = 32'b01111100000000000000000000000000;
                7'h46: rom_data = 32'b01111100000000000000000000000000;
                7'h47: rom_data = 32'b01111100000000000000000000000000;
                7'h48: rom_data = 32'b01111100000000000000000000000000;
                7'h49: rom_data = 32'b01111100000000000000000000000000; 
                7'h4A: rom_data = 32'b01111100000000000000000000000000;
                7'h4B: rom_data = 32'b01111100000000000000000000000000;
                7'h4C: rom_data = 32'b01111111111111111111111111111000;
                7'h4D: rom_data = 32'b01111111111111111111111111111000;
                7'h4E: rom_data = 32'b01111111111111111111111111111111;
                7'h4f: rom_data = 32'b01111111111111111111111111111111;
                7'h50: rom_data = 32'b01111111111111111111111111111111;
                7'h51: rom_data = 32'b00001111111111111111111111111111;
                7'h52: rom_data = 32'b00001111111111111111111111111111;
                7'h53: rom_data = 32'b00000000000000000000000001111111;
                7'h54: rom_data = 32'b00000000000000000000000001111111;
                7'h55: rom_data = 32'b00000000000000000000000001111111;
                7'h56: rom_data = 32'b00000000000000000000000001111111;
                7'h57: rom_data = 32'b00000000000000000000000001111111;
                7'h58: rom_data = 32'b00000000000000000000000001111111;
                7'h59: rom_data = 32'b01111111111111111111111111111111;
                7'h5a: rom_data = 32'b01111111111111111111111111111111;
                7'h5b: rom_data = 32'b01111111111111111111111111111111;
                7'h5c: rom_data = 32'b01111111111111111111111111111111;
                7'h5d: rom_data = 32'b01111111111111111111111111111000;
                7'h5e: rom_data = 32'b00011111111111111111111111111000;
                7'h5f: rom_data = 32'b00000000000000000000000000000000;
           endcase
endmodule